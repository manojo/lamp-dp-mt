-- VHDL Model Created for system "definition.vhd" 
-- 25/4/2010 18:25:36.277528
-- by Alpha2Vhdl Version 0.9 
