-- VHDL Model Created for system "definition.vhd" 
-- 5/1/2009 21:53:23.794258
-- by Alpha2Vhdl Version 0.9 
