-- VHDL Model Created for "system fir" 
-- 25/4/2010 18:24:33.427286
-- Alpha2Vhdl Version 0.9 
LIBRARY IEEE;
USE IEEE.std_logic_1164.all;
USE IEEE.std_logic_signed.all;
USE IEEE.numeric_std.all;

PACKAGE TYPES IS
  TYPE Array4To100OfInteger IS  ARRAY (4 TO 100) OF  SIGNED (15 DOWNTO 0);
END TYPES;

