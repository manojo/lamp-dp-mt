-- VHDL Model Created for system "definition.vhd" 
-- 23/4/2010 14:36:45.038174
-- by Alpha2Vhdl Version 0.9 
