-- VHDL Model Created for system "definition.vhd" 
-- 23/4/2010 8:38:34.239600
-- by Alpha2Vhdl Version 0.9 
