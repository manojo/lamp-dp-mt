-- VHDL Model Created for "system cellmatmultModule8" 
-- 29/12/2008 10:40:29.122989
-- Alpha2Vhdl Version 0.9 

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_signed.all;
use IEEE.numeric_std.all;

ENTITY cellmatmultModule8 IS
PORT(
  clk: IN STD_LOGIC;
  CE : IN STD_LOGIC;
  Rst : IN STD_LOGIC;
  C : OUT  SIGNED (15 DOWNTO 0)
);
END cellmatmultModule8;

ARCHITECTURE behavioural OF cellmatmultModule8 IS


  -- Insert missing components here!---------
   -- $MissingComponents$
BEGIN

    C <= "0000000000000000";

END behavioural;

