-- VHDL Model Created for "system computeDistances" 
-- 25/4/2010 18:25:37.044863
-- Alpha2Vhdl Version 0.9 
LIBRARY IEEE;
USE IEEE.std_logic_1164.all;
USE IEEE.std_logic_signed.all;
USE IEEE.numeric_std.all;

PACKAGE TYPES IS
  TYPE Array0To99OfSigned14To0 IS  ARRAY (0 TO 99) OF  SIGNED (14 DOWNTO 0);
END TYPES;

