-- VHDL Model Created for system "definition.vhd" 
-- 5/1/2009 21:53:46.231596
-- by Alpha2Vhdl Version 0.9 
