-- VHDL Model Created for system "definition.vhd" 
-- 23/4/2010 14:23:32.857114
-- by Alpha2Vhdl Version 0.9 
