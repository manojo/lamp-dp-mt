-- VHDL Model Created for system "definition.vhd" 
-- 23/4/2010 8:53:7.779618
-- by Alpha2Vhdl Version 0.9 
