-- VHDL Model Created for "system cellFirModule1" 
-- 15/7/2003 0:34:28
-- Alpha2Vhdl Version 0.9 

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_signed.all;
use IEEE.numeric_std.all;

ENTITY cellFirModule1 IS
PORT(
  Ck: IN STD_LOGIC;
  CE : IN STD_LOGIC;
  Rst : IN STD_LOGIC;
  H_mirr1 : IN  INTEGER RANGE -32768 TO 32767;
  x_mirr1 : IN  INTEGER RANGE -32768 TO 32767;
  Y : OUT  INTEGER RANGE -32768 TO 32767;
  xPipe : OUT  INTEGER RANGE -32768 TO 32767;
  HPipeES : OUT  INTEGER RANGE -32768 TO 32767;
  xPipeES : OUT  INTEGER RANGE -32768 TO 32767
);
END cellFirModule1;

ARCHITECTURE behavioural OF cellFirModule1 IS
    SIGNAL xPipeESloc4 :  INTEGER RANGE -32768 TO 32767 := 0;


  -- Insert missing components here!---------
BEGIN

    xPipeES <= xPipeESloc4;

    xPipeESloc4 <= x_mirr1;

    HPipeES <= H_mirr1;

    xPipe <= xPipeESloc4;

    Y <= 0;

END behavioural;

