library IEEE;
 use IEEE.std_logic_1164.all;
 Package definition is 

type B_In1Type is array (0 to 0) of Integer range -32767 to 32767;
type B_In_reg4locType is array (1 to 16) of Integer range -32767 to 32767;
type B_In2Type is array (1 to 15) of Integer range -32767 to 32767;
end definition; 

