-- VHDL Model Created for "system computeDistancesModule" 
-- 25/4/2010 18:25:36.904699
-- Alpha2Vhdl Version 0.9 
LIBRARY IEEE;
USE IEEE.std_logic_1164.all;
USE IEEE.std_logic_signed.all;
USE IEEE.numeric_std.all;

PACKAGE TYPES IS
  TYPE Array0To99OfBoolean IS  ARRAY (0 TO 99) OF  STD_LOGIC;
  TYPE Array0To99OfSigned14To0 IS  ARRAY (0 TO 99) OF  SIGNED (14 DOWNTO 0);
END TYPES;

