-- VHDL Model Created for system "definition.vhd" 
-- 25/4/2010 18:24:32.401029
-- by Alpha2Vhdl Version 0.9 
