library IEEE;
 use IEEE.std_logic_1164.all;
 Package definition is 

type Ilam1Type is array (1 to 1) of Integer range -32767 to 32767;
type Ilam2Type is array (1 to 1) of Integer range -32767 to 32767;
type Ix1Type is array (1 to 1) of Integer range -32767 to 32767;
type Ix2Type is array (1 to 1) of Integer range -32767 to 32767;
type Iy1Type is array (1 to 1) of Integer range -32767 to 32767;
type Iy2Type is array (1 to 1) of Integer range -32767 to 32767;
type Sl1Type is array (5 to 5) of Integer range -32767 to 32767;
type Sl2Type is array (5 to 5) of Integer range -32767 to 32767;
type SxType is array (5 to 5) of Integer range -32767 to 32767;
type SyType is array (5 to 5) of Integer range -32767 to 32767;
type Ol1Type is array (2 to 5) of Integer range -32767 to 32767;
type Ol2Type is array (2 to 5) of Integer range -32767 to 32767;
type OxType is array (2 to 5) of Integer range -32767 to 32767;
type OyType is array (2 to 5) of Integer range -32767 to 32767;
type OOl1Type is array (1 to 1) of Integer range -32767 to 32767;
type OOl2Type is array (1 to 1) of Integer range -32767 to 32767;
type OOxType is array (1 to 1) of Integer range -32767 to 32767;
type OOyType is array (1 to 1) of Integer range -32767 to 32767;
type IIl1Type is array (2 to 5) of Integer range -32767 to 32767;
type IIl2Type is array (2 to 5) of Integer range -32767 to 32767;
type IIxType is array (2 to 5) of Integer range -32767 to 32767;
type IIyType is array (2 to 5) of Integer range -32767 to 32767;
end definition; 

