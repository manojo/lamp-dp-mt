-- VHDL Model Created for "system firr" 
-- 23/4/2010 8:38:37.097264
-- Alpha2Vhdl Version 0.9 
LIBRARY IEEE;
USE IEEE.std_logic_1164.all;
USE IEEE.std_logic_signed.all;
USE IEEE.numeric_std.all;

PACKAGE TYPES IS
  TYPE Array-1To2OfInteger IS  ARRAY (-1 TO 2) OF  SIGNED (15 DOWNTO 0);
END TYPES;

