-- VHDL Model Created for system "definition.vhd" 
-- 5/1/2009 21:54:13.457973
-- by Alpha2Vhdl Version 0.9 
